module sbox (inp, outp);

input [3:0] inp;
output [3:0] outp;

reg [3:0] outp;

// implement the SBox design based on the truth table / boolean equations provided
// you can either use a high level concurrency construct or you can use continuous assignments


endmodule
